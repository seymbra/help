`timescale 1ns / 1ps
module xvga(input vclock_in,
            output reg [11:0] hcount_out,    // pixel number on current line
            output reg [10:0] vcount_out,     // line number
            output reg vsync_out, hsync_out,
            output reg blank_out);

   parameter DISPLAY_WIDTH  = 1024;      // display width
   parameter DISPLAY_HEIGHT = 768;       // number of lines

   parameter  H_FP = 24;                 // horizontal front porch
   parameter  H_SYNC_PULSE = 136;        // horizontal sync
   parameter  H_BP = 460;                // horizontal back porch

   parameter  V_FP = 3;                  // vertical front porch
   parameter  V_SYNC_PULSE = 6;          // vertical sync 
   parameter  V_BP = 29;                 // vertical back porch

   // horizontal: 1344 pixels total
   // display 1024 pixels per line
   reg hblank,vblank;
   wire hsyncon,hsyncoff,hreset,hblankon;
   assign hblankon = (hcount_out == (DISPLAY_WIDTH -1));    
   assign hsyncon = (hcount_out == (DISPLAY_WIDTH + H_FP - 1));  //1047
   assign hsyncoff = (hcount_out == (DISPLAY_WIDTH + H_FP + H_SYNC_PULSE - 1));  // 1183
   assign hreset = (hcount_out == (DISPLAY_WIDTH + H_FP + H_SYNC_PULSE + H_BP - 1));  //1343

   // vertical: 806 lines total
   // display 768 lines
   wire vsyncon,vsyncoff,vreset,vblankon;
   assign vblankon = hreset & (vcount_out == (DISPLAY_HEIGHT - 1));   // 767 
   assign vsyncon = hreset & (vcount_out == (DISPLAY_HEIGHT + V_FP - 1));  // 771
   assign vsyncoff = hreset & (vcount_out == (DISPLAY_HEIGHT + V_FP + V_SYNC_PULSE - 1));  // 777
   assign vreset = hreset & (vcount_out == (DISPLAY_HEIGHT + V_FP + V_SYNC_PULSE + V_BP - 1)); // 805

   // sync and blanking
   wire next_hblank,next_vblank;
   assign next_hblank = hreset ? 0 : hblankon ? 1 : hblank;
   assign next_vblank = vreset ? 0 : vblankon ? 1 : vblank;
   always_ff @(posedge vclock_in) begin
      hcount_out <= hreset ? 0 : hcount_out + 1;
      hblank <= next_hblank;
      hsync_out <= hsyncon ? 0 : hsyncoff ? 1 : hsync_out;  // active low

      vcount_out <= hreset ? (vreset ? 0 : vcount_out + 1) : vcount_out;
      vblank <= next_vblank;
      vsync_out <= vsyncon ? 0 : vsyncoff ? 1 : vsync_out;  // active low

      blank_out <= next_vblank | (next_hblank & ~hreset);
   end
   
endmodule


//`timescale 1ns / 1ps
//module xvga(input vclock_in,
//            output reg [10:0] hcount_out,    // pixel number on current line
//            output reg [9:0] vcount_out,     // line number
//            output reg vsync_out, hsync_out,
//            output reg blank_out);

//   parameter DISPLAY_WIDTH  = 1024;      // display width
//   parameter DISPLAY_HEIGHT = 768;       // number of lines

//   parameter  H_FP = 24;                 // horizontal front porch
//   parameter  H_SYNC_PULSE = 136;        // horizontal sync
//   parameter  H_BP = 160;                // horizontal back porch

//   parameter  V_FP = 3;                  // vertical front porch
//   parameter  V_SYNC_PULSE = 6;          // vertical sync 
//   parameter  V_BP = 29;                 // vertical back porch

//   // horizontal: 1344 pixels total
//   // display 1024 pixels per line
//   reg hblank,vblank;
//   wire hsyncon,hsyncoff,hreset,hblankon;
//   assign hblankon = (hcount_out == (DISPLAY_WIDTH -1));    
//   assign hsyncon = (hcount_out == (DISPLAY_WIDTH + H_FP - 1));  //1047
//   assign hsyncoff = (hcount_out == (DISPLAY_WIDTH + H_FP + H_SYNC_PULSE - 1));  // 1183
//   assign hreset = (hcount_out == (DISPLAY_WIDTH + H_FP + H_SYNC_PULSE + H_BP - 1));  //1343

//   // vertical: 806 lines total
//   // display 768 lines
//   wire vsyncon,vsyncoff,vreset,vblankon;
//   assign vblankon = hreset & (vcount_out == (DISPLAY_HEIGHT - 1));   // 767 
//   assign vsyncon = hreset & (vcount_out == (DISPLAY_HEIGHT + V_FP - 1));  // 771
//   assign vsyncoff = hreset & (vcount_out == (DISPLAY_HEIGHT + V_FP + V_SYNC_PULSE - 1));  // 777
//   assign vreset = hreset & (vcount_out == (DISPLAY_HEIGHT + V_FP + V_SYNC_PULSE + V_BP - 1)); // 805

//   // sync and blanking
//   wire next_hblank,next_vblank;
//   assign next_hblank = hreset ? 0 : hblankon ? 1 : hblank;
//   assign next_vblank = vreset ? 0 : vblankon ? 1 : vblank;
//   always_ff @(posedge vclock_in) begin
//      hcount_out <= hreset ? 0 : hcount_out + 1;
//      hblank <= next_hblank;
//      hsync_out <= hsyncon ? 0 : hsyncoff ? 1 : hsync_out;  // active low

//      vcount_out <= hreset ? (vreset ? 0 : vcount_out + 1) : vcount_out;
//      vblank <= next_vblank;
//      vsync_out <= vsyncon ? 0 : vsyncoff ? 1 : vsync_out;  // active low

//      blank_out <= next_vblank | (next_hblank & ~hreset);
//   end
   
//endmodule
